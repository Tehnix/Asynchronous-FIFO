package constants_pkg is
  constant DATA_WIDTH    : integer := 8;
  constant ADDRESS_WIDTH : integer := 5;
end constants_pkg;
